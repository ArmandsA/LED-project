-- Main entity

library ieee;
use ieee.std_logic_1164.all;

entity single_port_ram is



end entity;

architecture rtl of single_port_ram is

	
begin

	

end rtl;
